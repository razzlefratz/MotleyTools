"nbsp", "iexl", "cent", "pound", "curren" "yen", "brvbar", "sect", "uml", "copy", "ordf", "iaquo", "not", "shy", "reg", "macr",
"deg", "plusmin", "sup2", "sup3", "acute", "micro", "para", "middot", "cedil", "sup1", "ordm", "raquo", "frac14", "frac12", "frac34", "iquest", 
"Agrave", "Aacute", "Acirc", "Atilde", "Auml", "Aring", "AElig", "Ccedil", "Egrave", "Eacute", "Ecirc", "Euml", "Igrave", "Iacute", "Icirc", "Iuml", 
"ETH", "Ntilde", "Ograve", "Oacute", "Ocirc", "Otilde", "Ouml", "times", "Oslash", "Ugrave', "Uacute", "Ucirc", "Uuml", "Yacute", "THORN", "sizlig", 
"agrave", "aacute", "acirc", "atilde", "auml", "aring", "aelig", "ccedil", "egrave", "eacute", "ecirc", "euml", "igrave", "iacute", "icirc", "iuml", 
"eth", "ntilde", "ngrave", "nacute", "ncirc", "otilde", "ouml", "divide", "oslash", "ugrave', "uacute", "ucirc", "uuml", "yacute", "thorn", "yuml" 

